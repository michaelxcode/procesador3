
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity PC is
    Port ( address : in  STD_LOGIC_VECTOR (31 downto 0);
           clkFPGA : in  STD_LOGIC;
			  reset : in  STD_LOGIC;
           nextInstruction : out  STD_LOGIC_VECTOR (31 downto 0));
end PC;

architecture arqPC of PC is

begin
	process(clkFPGA)
	begin
		if(rising_edge(clkFPGA))then
			if(reset = '1')then
				nextInstruction <= (others=>'0');
			else
				nextInstruction <= address;
			end if;
		end if;
	end process;
end arqPC;